`include "src/misc_defines.header.sv"

//module Mux2To1(input logic a, b, sel,
//	output logic out);
//
//	always_comb
//	begin
//		out = (!sel) ? a : b;
//	end
//
//endmodule

module TestInstrDecoder;

	parameter __ARR_SIZE__MAX_NUM_INSTRUCTIONS = 1024;
	parameter __LAST_INDEX__MAX_NUM_INSTRUCTIONS 
		= `ARR_SIZE_TO_LAST_INDEX(__ARR_SIZE__MAX_NUM_INSTRUCTIONS);

	logic [`MSB_POS__INSTRUCTION:0] 
		__instructions[0 : __LAST_INDEX__MAX_NUM_INSTRUCTIONS];

	initial
	begin
		$readmemh("instructions.txt.ignore", __instructions);
	end



	// Stuffs!
endmodule
