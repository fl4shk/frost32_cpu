`ifndef src__slash__main_mem_defines_header_sv
`define src__slash__main_mem_defines_header_sv

// src/main_mem_defines.header.sv

`include "src/misc_defines.header.sv"

//`define WIDTH__MAIN_MEM_

`endif		// src__slash__main_mem_defines_header_sv
