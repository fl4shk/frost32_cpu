`ifndef src__slash__instr_decoder_stuff_header_sv
`define src__slash__instr_decoder_stuff_header_sv

// src/instr_decoder_stuff.header.sv

`include "src/misc_defines.header.sv"

`define INSTR_DEC__WIDTH_OP 4
`define INSTR_DEC__MSB_POS_OP `WIDTH_TO_MSB_POS(`INSTR_DEC__WIDTH_OP)

`endif		// src__slash__instr_decoder_stuff_header_sv
