`include "src/instr_decoder_defines.header.sv"


