`include "src/cache_defines.header.sv"
