module TopLevel;
	
endmodule
